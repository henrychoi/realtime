module application#(parameter DELAY=1, SYNC_WINDOW=1, FP_SIZE=1, N_PATCH=1
, N_CAM=1)
( input CLK, RESET, output[7:0] GPIO_LED);
`include "function.v"
endmodule
